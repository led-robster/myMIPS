


module top #(
    parameters
) (
    
);







    
endmodule