

// module btt_generator #(
//     parameters
// ) (
//     ports
// );
    
// endmodule